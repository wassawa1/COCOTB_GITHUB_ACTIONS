module dff (
    input wire clk,
    input wire reset,
    input wire d,
    output reg q
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        q <= 0;  // Reset value
    end else begin
        q <= d;
    end
end

endmodule
